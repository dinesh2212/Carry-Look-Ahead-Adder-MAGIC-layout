magic
tech scmos
timestamp 1619620769
<< nwell >>
rect -43 -14 9 22
rect 53 -14 94 23
rect 169 -9 221 27
<< ntransistor >>
rect 73 -39 75 -29
rect -23 -64 -21 -54
rect -9 -64 -7 -54
rect 189 -59 191 -49
rect 203 -59 205 -49
<< ptransistor >>
rect -23 -6 -21 14
rect -9 -6 -7 14
rect 73 -6 75 14
rect 189 -1 191 19
rect 203 -1 205 19
<< ndiffusion >>
rect 69 -39 73 -29
rect 75 -39 79 -29
rect -27 -64 -23 -54
rect -21 -64 -9 -54
rect -7 -64 -3 -54
rect 185 -59 189 -49
rect 191 -59 203 -49
rect 205 -59 209 -49
<< pdiffusion >>
rect -27 -6 -23 14
rect -21 -6 -9 14
rect -7 -6 -3 14
rect 69 -6 73 14
rect 75 -6 79 14
rect 185 -1 189 19
rect 191 -1 203 19
rect 205 -1 209 19
<< ndcontact >>
rect 65 -39 69 -29
rect 79 -39 83 -29
rect -31 -64 -27 -54
rect -3 -64 1 -54
rect 181 -59 185 -49
rect 209 -59 213 -49
<< pdcontact >>
rect -31 -6 -27 14
rect -3 -6 1 14
rect 65 -6 69 14
rect 79 -6 83 14
rect 181 -1 185 19
rect 209 -1 213 19
<< polysilicon >>
rect -23 14 -21 17
rect -9 14 -7 17
rect 73 14 75 17
rect 110 16 112 59
rect 124 24 154 26
rect 189 19 191 22
rect 203 19 205 22
rect -23 -54 -21 -6
rect -9 -25 -7 -6
rect 73 -29 75 -6
rect 143 -18 145 6
rect -9 -54 -7 -33
rect 73 -42 75 -39
rect 161 -42 163 -16
rect 189 -49 191 -1
rect 203 -20 205 -1
rect 203 -49 205 -28
rect 189 -62 191 -59
rect 203 -62 205 -59
rect -23 -67 -21 -64
rect -9 -67 -7 -64
rect 31 -115 33 -73
rect 121 -74 150 -72
<< polycontact >>
rect 112 55 116 59
rect 120 23 124 27
rect 150 26 154 30
rect 109 12 113 16
rect 142 6 146 10
rect -27 -15 -23 -11
rect -13 -25 -9 -21
rect 69 -23 73 -19
rect 185 -10 189 -6
rect 142 -22 146 -18
rect -13 -37 -9 -33
rect 163 -20 167 -16
rect 160 -46 164 -42
rect 199 -20 203 -16
rect 199 -32 203 -28
rect 30 -73 34 -69
rect 117 -75 121 -71
rect 150 -75 154 -71
rect 33 -115 37 -111
<< metal1 >>
rect 116 55 145 59
rect -71 45 -66 46
rect -71 41 146 45
rect -71 -21 -66 41
rect -46 23 120 27
rect -31 14 -27 23
rect 65 14 69 23
rect -54 -15 -27 -11
rect -79 -25 -13 -21
rect -79 -37 -13 -33
rect -73 -88 -69 -37
rect -3 -45 1 -6
rect 79 -18 83 -6
rect 109 -6 113 12
rect 142 10 146 41
rect 150 30 232 32
rect 154 28 232 30
rect 181 19 185 28
rect 109 -10 185 -6
rect 109 -18 113 -10
rect 21 -23 69 -19
rect 79 -22 113 -18
rect 167 -20 199 -16
rect 21 -45 26 -23
rect -31 -49 26 -45
rect -3 -54 1 -49
rect -31 -76 -27 -64
rect 30 -69 34 -23
rect 79 -29 83 -22
rect 142 -28 146 -22
rect 142 -32 199 -28
rect 65 -45 69 -39
rect 209 -40 213 -1
rect 53 -49 98 -45
rect 181 -44 251 -40
rect 61 -71 65 -49
rect 131 -50 164 -46
rect 209 -49 213 -44
rect 61 -75 117 -71
rect 61 -76 65 -75
rect -49 -80 65 -76
rect 131 -88 135 -50
rect 181 -71 185 -59
rect 154 -75 229 -71
rect -73 -92 135 -88
rect 247 -111 251 -44
rect 37 -115 251 -111
<< labels >>
rlabel metal1 -46 23 120 27 1 vdd
rlabel metal1 53 -49 98 -45 1 gnd
rlabel metal1 -54 -15 -27 -11 1 in_D
rlabel metal1 -79 -25 -13 -21 1 in_en_bar
rlabel metal1 -79 -37 -13 -33 1 in_en
rlabel metal1 83 -22 113 -18 1 q_out
<< end >>
