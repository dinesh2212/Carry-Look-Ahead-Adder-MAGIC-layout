magic
tech scmos
timestamp 1618919255
<< polysilicon >>
rect 107 88 140 90
<< polycontact >>
rect 136 90 140 94
rect 107 84 111 88
<< metal1 >>
rect -36 331 130 335
rect -36 174 -32 331
rect -149 170 -102 174
rect -68 170 -21 174
rect -135 125 -131 170
rect -25 132 -21 170
rect -25 128 0 132
rect -135 121 0 125
rect 126 121 130 331
rect -135 114 0 118
rect 126 117 149 121
rect -135 47 -131 114
rect -25 107 0 111
rect 136 110 149 114
rect -25 47 -21 107
rect 93 95 125 99
rect -149 43 -102 47
rect -68 43 -21 47
rect -39 -11 -35 43
rect 107 -11 111 84
rect 121 71 125 95
rect 136 94 140 110
rect 194 103 224 107
rect 121 67 224 71
rect -39 -15 111 -11
use inv_2W  inv_2W_0
timestamp 1618844995
transform 1 0 -81 0 1 183
box -21 -45 13 49
use inv_2W  inv_2W_1
timestamp 1618844995
transform 1 0 -81 0 1 56
box -21 -45 13 49
use xor_4W  xor_4W_0
timestamp 1618844952
transform 1 0 37 0 1 151
box -37 -151 56 172
use and  and_0
timestamp 1618746604
transform 1 0 180 0 1 127
box -31 -48 16 55
<< end >>
