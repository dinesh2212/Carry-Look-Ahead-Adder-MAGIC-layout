magic
tech scmos
timestamp 1619594738
<< polysilicon >>
rect -9 1643 26 1645
rect 30 1560 32 1583
rect -63 1422 -9 1424
rect -22 1406 29 1408
rect -6 1387 33 1389
rect -32 1374 10 1376
rect -79 1353 -13 1355
rect -98 1332 -9 1334
<< polycontact >>
rect -9 1639 -5 1643
rect 26 1642 30 1646
rect 29 1583 33 1587
rect 29 1556 33 1560
rect -63 1418 -59 1422
rect -9 1421 -5 1425
rect -26 1405 -22 1409
rect 29 1405 33 1409
rect 29 1389 33 1393
rect -6 1383 -2 1387
rect -32 1370 -28 1374
rect 10 1373 14 1377
rect -79 1349 -75 1353
rect -13 1352 -9 1356
rect -13 1334 -9 1338
rect -98 1328 -94 1332
<< metal1 >>
rect 10 1650 50 1654
rect -9 1425 -5 1639
rect -98 475 -94 1328
rect -79 488 -75 1349
rect -63 500 -59 1418
rect -48 1405 -26 1409
rect -48 512 -44 1405
rect -9 1400 -5 1421
rect -15 1396 -5 1400
rect -32 523 -28 1370
rect -15 1363 -11 1396
rect -6 1370 -2 1383
rect 10 1377 14 1650
rect 30 1642 50 1646
rect 29 1634 58 1638
rect 29 1587 33 1634
rect 29 1409 33 1556
rect 29 1393 33 1405
rect 14 1373 39 1377
rect -6 1366 39 1370
rect -15 1359 39 1363
rect -9 1352 39 1356
rect -13 1345 39 1349
rect -13 1338 -9 1345
rect -32 519 8 523
rect -48 508 8 512
rect -63 496 8 500
rect -79 484 8 488
rect -98 471 8 475
rect -106 460 8 464
rect -106 449 8 453
use c2  c2_0
timestamp 1619090282
transform 1 0 89 0 1 1662
box -39 -78 46 56
use c3  c3_0
timestamp 1619526073
transform 1 0 106 0 1 1389
box -78 -171 55 185
use c4  c4_0
timestamp 1619545755
transform 1 0 75 0 1 541
box -75 -541 152 662
<< end >>
