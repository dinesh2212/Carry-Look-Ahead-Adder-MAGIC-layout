magic
tech scmos
timestamp 1618898111
<< nwell >>
rect -22 -15 46 77
<< ntransistor >>
rect -10 -100 -8 -60
rect 4 -100 6 -60
rect 18 -100 20 -60
rect 32 -100 34 -60
<< ptransistor >>
rect -10 -9 -8 71
rect 4 -9 6 71
rect 18 -9 20 71
rect 32 -9 34 71
<< ndiffusion >>
rect -12 -100 -10 -60
rect -8 -100 4 -60
rect 6 -100 10 -60
rect 14 -100 18 -60
rect 20 -100 32 -60
rect 34 -100 36 -60
<< pdiffusion >>
rect -12 -9 -10 71
rect -8 -9 -4 71
rect 0 -9 4 71
rect 6 -9 10 71
rect 14 -9 18 71
rect 20 -9 24 71
rect 28 -9 32 71
rect 34 -9 36 71
<< ndcontact >>
rect -16 -100 -12 -60
rect 10 -100 14 -60
rect 36 -100 40 -60
<< pdcontact >>
rect -16 -9 -12 71
rect -4 -9 0 71
rect 10 -9 14 71
rect 24 -9 28 71
rect 36 -9 40 71
<< polysilicon >>
rect -10 71 -8 74
rect 4 71 6 74
rect 18 71 20 74
rect 32 71 34 74
rect -10 -60 -8 -9
rect 4 -60 6 -9
rect 18 -60 20 -9
rect 32 -60 34 -9
rect -10 -103 -8 -100
rect 4 -103 6 -100
rect 18 -103 20 -100
rect 32 -103 34 -100
<< polycontact >>
rect -14 -33 -10 -29
rect 0 -40 4 -36
rect 14 -47 18 -43
rect 28 -26 32 -22
<< metal1 >>
rect -27 85 51 89
rect -4 71 0 85
rect 10 77 40 81
rect 10 71 14 77
rect 36 71 40 77
rect -16 -15 -12 -9
rect 10 -15 14 -9
rect -16 -19 14 -15
rect 24 -15 28 -9
rect 24 -19 48 -15
rect -34 -26 28 -22
rect -34 -33 -14 -29
rect -34 -40 0 -36
rect -34 -47 14 -43
rect 44 -51 48 -19
rect -16 -55 51 -51
rect -16 -60 -12 -55
rect 36 -60 40 -55
rect 10 -107 14 -100
rect -27 -111 51 -107
<< labels >>
rlabel metal1 -27 -111 51 -107 1 gnd
rlabel metal1 -27 85 51 89 5 vdd
rlabel metal1 -16 -55 51 -51 1 out
rlabel metal1 -34 -26 28 -22 1 in_a_bar
rlabel metal1 -34 -33 -14 -29 1 in_a
rlabel metal1 -34 -40 0 -36 1 in_b
rlabel metal1 -34 -47 14 -43 1 in_b_bar
<< end >>
