magic
tech scmos
timestamp 1618746604
<< nwell >>
rect -25 -8 11 52
<< ntransistor >>
rect -13 -39 -11 -27
rect -3 -39 -1 -27
<< ptransistor >>
rect -13 -2 -11 46
rect -3 -2 -1 46
<< ndiffusion >>
rect -15 -39 -13 -27
rect -11 -39 -9 -27
rect -5 -39 -3 -27
rect -1 -39 1 -27
<< pdiffusion >>
rect -15 -2 -13 46
rect -11 -2 -3 46
rect -1 -2 1 46
<< ndcontact >>
rect -19 -39 -15 -27
rect -9 -39 -5 -27
rect 1 -39 5 -27
<< pdcontact >>
rect -19 -2 -15 46
rect 1 -2 5 46
<< polysilicon >>
rect -13 46 -11 49
rect -3 46 -1 49
rect -13 -27 -11 -2
rect -3 -27 -1 -2
rect -13 -42 -11 -39
rect -3 -42 -1 -39
<< polycontact >>
rect -17 -10 -13 -6
rect -7 -17 -3 -13
<< metal1 >>
rect -30 51 16 55
rect -19 46 -15 51
rect -31 -10 -17 -6
rect -31 -17 -7 -13
rect 1 -20 5 -2
rect -19 -24 14 -20
rect -9 -27 -5 -24
rect -19 -44 -15 -39
rect 1 -44 5 -39
rect -30 -48 16 -44
<< labels >>
rlabel metal1 -31 -10 -17 -6 1 in1
rlabel metal1 -31 -17 -7 -13 1 in2
rlabel metal1 -19 -24 14 -20 1 out
rlabel metal1 -30 51 16 55 5 vdd
rlabel metal1 -30 -48 16 -44 1 gnd
<< end >>
