magic
tech scmos
timestamp 1619631775
<< polysilicon >>
rect 1771 2119 1800 2121
rect 1789 1747 1819 1749
rect 479 1595 481 1632
rect 574 1586 576 1674
rect 608 1586 610 1661
rect 1193 1618 1195 1647
rect 1350 1583 1352 1674
rect 1376 1583 1378 1661
rect 1097 1418 1137 1420
rect 1790 1413 1819 1415
rect 1399 1193 1401 1216
rect 354 1049 356 1076
rect 380 1051 382 1079
rect 479 1038 481 1085
rect 574 1047 576 1082
rect 608 1047 610 1082
rect 1781 1080 1814 1082
rect 653 1062 746 1064
rect 380 832 382 860
rect -9 801 -7 827
rect 574 650 576 681
rect 608 650 610 681
rect 653 660 730 662
rect 574 578 576 615
rect 608 576 610 619
rect 653 596 715 598
rect 393 418 395 447
rect 608 409 610 453
rect 659 430 699 432
rect 1246 299 1312 301
rect 1785 293 1814 295
rect 1264 -209 1266 -173
<< polycontact >>
rect 1767 2118 1771 2122
rect 1800 2118 1804 2122
rect 1785 1746 1789 1750
rect 1819 1746 1823 1750
rect 481 1628 485 1632
rect 478 1591 482 1595
rect 576 1670 580 1674
rect 1346 1670 1350 1674
rect 610 1657 614 1661
rect 1189 1643 1193 1647
rect 1195 1618 1199 1622
rect 573 1582 577 1586
rect 607 1582 611 1586
rect 1372 1657 1376 1661
rect 1349 1579 1353 1583
rect 1375 1579 1379 1583
rect 1093 1417 1097 1421
rect 1137 1417 1141 1421
rect 1786 1412 1790 1416
rect 1819 1412 1823 1416
rect 1398 1216 1402 1220
rect 1401 1193 1405 1197
rect 478 1085 482 1089
rect 353 1076 357 1080
rect 379 1079 383 1083
rect 353 1045 357 1049
rect 379 1047 383 1051
rect 573 1082 577 1086
rect 607 1082 611 1086
rect 1777 1079 1781 1083
rect 1814 1079 1818 1083
rect 649 1061 653 1065
rect 746 1061 750 1065
rect 573 1043 577 1047
rect 607 1043 611 1047
rect 478 1034 482 1038
rect 379 860 383 864
rect -10 827 -6 831
rect 379 828 383 832
rect -10 797 -6 801
rect 573 681 577 685
rect 607 681 611 685
rect 649 659 653 663
rect 730 659 734 663
rect 573 646 577 650
rect 607 646 611 650
rect 607 619 611 623
rect 573 615 577 619
rect 573 574 577 578
rect 649 595 653 599
rect 715 595 719 599
rect 607 572 611 576
rect 607 453 611 457
rect 392 447 396 451
rect 392 414 396 418
rect 655 429 659 433
rect 699 429 703 433
rect 607 405 611 409
rect 1241 298 1246 302
rect 1312 298 1317 302
rect 1781 292 1785 296
rect 1814 292 1818 296
rect 1263 -173 1267 -169
rect 1263 -213 1267 -209
<< metal1 >>
rect 353 2155 358 2158
rect 353 2151 1732 2155
rect 353 1704 358 2151
rect 1728 2122 1732 2151
rect 1728 2118 1767 2122
rect 1701 1746 1785 1750
rect -996 1287 -988 1294
rect -996 1283 -22 1287
rect -996 1206 -988 1283
rect -1133 1199 -988 1206
rect -155 1205 -55 1209
rect -59 1049 -55 1205
rect -26 1139 -22 1283
rect -26 1135 20 1139
rect 353 1080 357 1704
rect 580 1670 1346 1674
rect 614 1657 1372 1661
rect 379 1643 1189 1647
rect 379 1083 383 1643
rect 485 1628 1432 1632
rect 1428 1624 1432 1628
rect 1199 1618 1407 1622
rect 1403 1617 1407 1618
rect 401 1611 1152 1615
rect 1403 1613 1428 1617
rect 401 1065 405 1611
rect 1148 1610 1152 1611
rect 1148 1606 1428 1610
rect 1399 1601 1428 1603
rect 521 1599 1428 1601
rect 521 1597 1402 1599
rect 478 1089 482 1591
rect 521 1065 525 1597
rect 1701 1595 1705 1746
rect 1564 1591 1705 1595
rect 573 1086 577 1582
rect 607 1086 611 1582
rect 913 1490 1032 1494
rect 1066 1490 1119 1494
rect 984 1421 988 1490
rect 984 1417 1093 1421
rect 1115 1392 1119 1490
rect 1141 1417 1325 1421
rect 1321 1399 1325 1417
rect 1349 1406 1353 1579
rect 1375 1413 1379 1579
rect 1375 1409 1427 1413
rect 1729 1412 1786 1416
rect 1349 1402 1427 1406
rect 1321 1395 1427 1399
rect 1115 1388 1427 1392
rect 1729 1384 1733 1412
rect 1563 1380 1733 1384
rect 1029 1255 1402 1259
rect 1029 1203 1033 1255
rect 1398 1220 1402 1255
rect 1359 1203 1427 1204
rect 939 1199 1055 1203
rect 1089 1200 1427 1203
rect 1089 1199 1363 1200
rect 1405 1193 1427 1197
rect 1263 1186 1427 1190
rect 369 1061 412 1065
rect 446 1061 649 1065
rect 369 1058 373 1061
rect -59 1045 20 1049
rect 353 1022 357 1045
rect -91 905 -87 906
rect -91 901 20 905
rect -868 897 -864 901
rect -91 897 -87 901
rect -868 891 -87 897
rect -868 847 -864 891
rect -1178 843 -863 847
rect -160 834 -34 838
rect -38 815 -34 834
rect -10 831 -6 901
rect 379 864 383 1047
rect 478 876 482 1034
rect 478 872 516 876
rect 368 844 416 848
rect 450 844 451 848
rect 368 824 372 844
rect -38 811 20 815
rect -38 618 -34 811
rect -10 693 -6 797
rect 368 768 372 786
rect 379 768 383 828
rect 512 768 516 872
rect 368 764 416 768
rect 450 764 516 768
rect -10 689 39 693
rect 573 685 577 1043
rect 607 685 611 1043
rect 352 659 415 663
rect 449 659 649 663
rect 352 650 356 659
rect 344 646 356 650
rect 573 619 577 646
rect 607 623 611 646
rect -38 614 39 618
rect 344 605 356 609
rect 352 599 356 605
rect 352 595 415 599
rect 449 595 649 599
rect -906 550 -902 553
rect -906 546 -48 550
rect -906 499 -902 546
rect -1157 495 -902 499
rect -52 498 -48 546
rect -52 494 21 498
rect -151 485 -88 490
rect 573 486 577 574
rect -92 408 -88 485
rect 392 482 577 486
rect 392 451 396 482
rect 607 457 611 572
rect 369 429 415 433
rect 449 429 655 433
rect 369 417 373 429
rect -92 404 21 408
rect 369 360 373 378
rect 392 360 396 414
rect 607 360 611 405
rect 369 356 415 360
rect 449 356 683 360
rect 483 323 672 327
rect -828 205 -75 206
rect -832 201 -75 205
rect -832 160 -828 201
rect -79 189 -75 201
rect -79 185 0 189
rect -1172 156 -828 160
rect -156 152 -96 156
rect -101 62 -97 152
rect 483 131 487 323
rect 369 127 415 131
rect 449 127 487 131
rect 523 312 672 316
rect 369 118 373 127
rect -101 58 0 62
rect 369 39 373 82
rect 523 39 527 312
rect 1005 298 1241 302
rect 369 35 415 39
rect 449 35 527 39
rect 381 -228 388 35
rect 495 -188 499 35
rect 1263 -169 1267 1186
rect 1294 1179 1427 1183
rect 1294 -188 1298 1179
rect 1563 1171 1706 1175
rect 1702 1083 1706 1171
rect 1702 1079 1777 1083
rect 1702 1078 1706 1079
rect 1317 298 1756 302
rect 1752 296 1756 298
rect 1752 292 1781 296
rect 495 -192 1298 -188
rect 1263 -228 1267 -213
rect 381 -232 1267 -228
use dflipflop  dflipflop_12
timestamp 1619621930
transform 1 0 1775 0 1 2018
box 0 -22 750 207
use dflipflop  dflipflop_4
timestamp 1619621930
transform 1 0 -1883 0 1 1031
box 0 -22 750 207
use dflipflop  dflipflop_0
timestamp 1619621930
transform 1 0 -905 0 1 1035
box 0 -22 750 207
use dflipflop  dflipflop_5
timestamp 1619621930
transform 1 0 -1903 0 1 673
box 0 -22 750 207
use dflipflop  dflipflop_1
timestamp 1619621930
transform 1 0 -910 0 1 664
box 0 -22 750 207
use dflipflop  dflipflop_6
timestamp 1619621930
transform 1 0 -1907 0 1 325
box 0 -22 750 207
use dflipflop  dflipflop_2
timestamp 1619621930
transform 1 0 -901 0 1 316
box 0 -22 750 207
use dflipflop  dflipflop_7
timestamp 1619621930
transform 1 0 -1922 0 1 -14
box 0 -22 750 207
use dflipflop  dflipflop_3
timestamp 1619621930
transform 1 0 -906 0 1 -18
box 0 -22 750 207
use pg  pg_0
timestamp 1618920172
transform 1 0 20 0 1 1002
box -20 -1002 353 220
use inv_W  inv_W_0
timestamp 1618656596
transform 1 0 427 0 1 1070
box -15 -30 19 31
use inv_W  inv_W_1
timestamp 1618656596
transform 1 0 431 0 1 853
box -15 -30 19 31
use inv_W  inv_W_2
timestamp 1618656596
transform 1 0 431 0 1 773
box -15 -30 19 31
use inv_W  inv_W_3
timestamp 1618656596
transform 1 0 430 0 1 668
box -15 -30 19 31
use inv_W_2  inv_W_2_0
timestamp 1618743374
transform 1 0 432 0 1 617
box -17 -39 17 10
use inv_W  inv_W_4
timestamp 1618656596
transform 1 0 430 0 1 438
box -15 -30 19 31
use inv_W  inv_W_5
timestamp 1618656596
transform 1 0 430 0 1 365
box -15 -30 19 31
use inv_W  inv_W_6
timestamp 1618656596
transform 1 0 430 0 1 136
box -15 -30 19 31
use inv_2W  inv_2W_0
timestamp 1618844995
transform 1 0 436 0 1 48
box -21 -45 13 49
use CLA  CLA_0
timestamp 1619594738
transform 1 0 778 0 1 -137
box -106 0 227 1718
use inv_W  inv_W_8
timestamp 1618656596
transform 1 0 1047 0 1 1499
box -15 -30 19 31
use inv_W  inv_W_7
timestamp 1618656596
transform 1 0 1070 0 1 1208
box -15 -30 19 31
use sum  sum_0
timestamp 1619597960
transform 1 0 1428 0 1 1535
box -1 -420 136 200
use dflipflop  dflipflop_8
timestamp 1619621930
transform 1 0 1794 0 1 1646
box 0 -22 750 207
use dflipflop  dflipflop_9
timestamp 1619621930
transform 1 0 1794 0 1 1312
box 0 -22 750 207
use dflipflop  dflipflop_10
timestamp 1619621930
transform 1 0 1789 0 1 979
box 0 -22 750 207
use dflipflop  dflipflop_11
timestamp 1619621930
transform 1 0 1789 0 1 192
box 0 -22 750 207
<< end >>
