magic
tech scmos
timestamp 1619090282
<< nwell >>
rect -30 -1 29 52
<< ntransistor >>
rect -16 -61 -14 -41
rect -2 -61 0 -41
rect 12 -61 14 -41
<< ptransistor >>
rect -16 5 -14 45
rect -2 5 0 45
rect 12 14 14 34
<< ndiffusion >>
rect -20 -61 -16 -41
rect -14 -61 -10 -41
rect -6 -61 -2 -41
rect 0 -61 4 -41
rect 8 -61 12 -41
rect 14 -61 18 -41
<< pdiffusion >>
rect -20 5 -16 45
rect -14 5 -2 45
rect 0 5 4 45
rect 8 14 12 34
rect 14 14 18 34
<< ndcontact >>
rect -24 -61 -20 -41
rect -10 -61 -6 -41
rect 4 -61 8 -41
rect 18 -61 22 -41
<< pdcontact >>
rect -24 5 -20 45
rect 4 14 8 34
rect 18 14 22 34
<< polysilicon >>
rect -16 45 -14 48
rect -2 45 0 48
rect 12 34 14 37
rect -16 -41 -14 5
rect -2 -41 0 5
rect 12 -41 14 14
rect -16 -64 -14 -61
rect -2 -64 0 -61
rect 12 -64 14 -61
<< polycontact >>
rect -20 -12 -16 -8
rect -6 -20 -2 -16
rect 8 -28 12 -24
<< metal1 >>
rect -38 52 37 56
rect 4 34 8 52
rect -24 1 -20 5
rect 18 1 22 14
rect -24 -3 27 1
rect -39 -12 -20 -8
rect -39 -20 -6 -16
rect -39 -28 8 -24
rect 23 -31 27 -3
rect -10 -35 46 -31
rect -10 -41 -6 -35
rect -24 -65 -20 -61
rect 4 -65 8 -61
rect -24 -69 8 -65
rect 18 -74 22 -61
rect -38 -78 37 -74
<< labels >>
rlabel metal1 -38 -78 37 -74 1 gnd
rlabel metal1 -38 52 37 56 5 vdd
rlabel metal1 -39 -12 -20 -8 1 in_g0_bar
rlabel metal1 -39 -20 -6 -16 1 in_p1_bar
rlabel metal1 -39 -28 8 -24 1 in_g1_bar
rlabel metal1 -10 -35 46 -31 1 c2_out
<< end >>
