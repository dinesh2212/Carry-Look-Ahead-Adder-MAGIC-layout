magic
tech scmos
timestamp 1619545755
<< nwell >>
rect -67 -12 113 655
<< ntransistor >>
rect -49 -398 -47 -318
rect -26 -438 -24 -278
rect -6 -398 -4 -318
rect 16 -438 18 -278
rect 38 -518 40 -198
rect 60 -518 62 -198
rect 82 -518 84 -198
<< ptransistor >>
rect -49 240 -47 400
rect -26 240 -24 400
rect -6 240 -4 400
rect 16 160 18 480
rect 38 160 40 480
rect 60 0 62 640
rect 82 0 84 640
<< ndiffusion >>
rect -53 -398 -49 -318
rect -47 -398 -34 -318
rect -30 -438 -26 -278
rect -24 -438 -22 -278
rect -10 -398 -6 -318
rect -4 -398 8 -318
rect 12 -438 16 -278
rect 18 -438 30 -278
rect 34 -518 38 -198
rect 40 -518 52 -198
rect 56 -518 60 -198
rect 62 -518 74 -198
rect 78 -518 82 -198
rect 84 -518 88 -198
<< pdiffusion >>
rect -52 240 -49 400
rect -47 240 -34 400
rect -30 240 -26 400
rect -24 240 -14 400
rect -10 240 -6 400
rect -4 240 0 400
rect 12 160 16 480
rect 18 160 30 480
rect 34 160 38 480
rect 40 160 52 480
rect 56 0 60 640
rect 62 0 82 640
rect 84 0 88 640
<< ndcontact >>
rect -57 -398 -53 -318
rect -34 -438 -30 -278
rect -22 -438 -18 -278
rect -14 -398 -10 -318
rect 8 -438 12 -278
rect 30 -518 34 -198
rect 52 -518 56 -198
rect 74 -518 78 -198
rect 88 -518 92 -198
<< pdcontact >>
rect -56 240 -52 400
rect -34 240 -30 400
rect -14 240 -10 400
rect 0 240 4 400
rect 8 160 12 480
rect 30 160 34 480
rect 52 0 56 640
rect 88 0 92 640
<< polysilicon >>
rect 60 640 62 643
rect 82 640 84 643
rect -49 400 -47 460
rect -26 400 -24 478
rect -6 400 -4 494
rect 16 480 18 483
rect 38 480 40 483
rect -49 -318 -47 240
rect -26 -278 -24 240
rect -49 -402 -47 -398
rect -6 -318 -4 240
rect 16 -278 18 160
rect 38 -198 40 160
rect 60 -198 62 0
rect 82 -198 84 0
rect -6 -402 -4 -398
rect -26 -442 -24 -438
rect 16 -442 18 -438
rect 38 -521 40 -518
rect 60 -521 62 -518
rect 82 -521 84 -518
<< polycontact >>
rect -53 -81 -49 -77
rect -30 -57 -26 -53
rect -10 -92 -6 -88
rect 12 -70 16 -66
rect 34 -33 38 -29
rect 56 -22 60 -18
rect 78 -45 82 -41
<< metal1 >>
rect -68 658 113 662
rect 0 411 4 658
rect 30 646 92 650
rect 30 480 34 646
rect 88 640 92 646
rect -56 407 4 411
rect -56 400 -52 407
rect 0 400 4 407
rect -34 -6 -30 240
rect -14 154 -10 240
rect 8 154 12 160
rect -14 150 12 154
rect 52 -6 56 0
rect -34 -7 56 -6
rect -34 -11 125 -7
rect -67 -22 56 -18
rect -67 -33 34 -29
rect -67 -45 78 -41
rect -67 -57 -30 -53
rect -67 -70 12 -66
rect -67 -81 -53 -77
rect -67 -92 -10 -88
rect 121 -102 125 -11
rect 121 -106 152 -102
rect 121 -191 125 -106
rect 8 -195 125 -191
rect -34 -273 -10 -269
rect -34 -278 -30 -273
rect -57 -537 -53 -398
rect -14 -318 -10 -273
rect 8 -278 12 -195
rect 74 -198 78 -195
rect -22 -526 -18 -438
rect 30 -526 34 -518
rect -22 -530 34 -526
rect 52 -526 56 -518
rect 88 -526 92 -518
rect 52 -530 92 -526
rect -75 -541 117 -537
<< labels >>
rlabel metal1 -68 658 113 662 5 vdd
rlabel metal1 -75 -541 117 -537 1 gnd
rlabel metal1 121 -106 152 -102 1 c4_out
rlabel metal1 -67 -22 56 -18 1 in_g0_bar
rlabel metal1 -67 -33 34 -29 1 in_g1_bar
rlabel metal1 -67 -45 78 -41 1 in_p1_bar
rlabel metal1 -67 -57 -30 -53 1 in_g2_bar
rlabel metal1 -67 -70 12 -66 1 in_p2_bar
rlabel metal1 -67 -81 -53 -77 1 in_g3_bar
rlabel metal1 -67 -92 -10 -88 1 in_p3_bar
<< end >>
